library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package emulate_bitstream is
--X0Y1, W_IO
constant Tile_X0Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011000000000000000011000001100000000000000000000000";
--X1Y1, LUT4AB
constant Tile_X1Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X2Y1, LUT4AB
constant Tile_X2Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X3Y1, RegFile
constant Tile_X3Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y1, LUT4AB
constant Tile_X4Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X5Y1, LUT4AB
constant Tile_X5Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000010000";
--X6Y1, DSP_top
constant Tile_X6Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y1, LUT4AB
constant Tile_X7Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X8Y1, LUT4AB
constant Tile_X8Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X9Y1, RAM_IO
constant Tile_X9Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y2, W_IO
constant Tile_X0Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000110000000000000000000000000011101111100000000000000000000000";
--X1Y2, LUT4AB
constant Tile_X1Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000";
--X2Y2, LUT4AB
constant Tile_X2Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X3Y2, RegFile
constant Tile_X3Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y2, LUT4AB
constant Tile_X4Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X5Y2, LUT4AB
constant Tile_X5Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X6Y2, DSP_bot
constant Tile_X6Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y2, LUT4AB
constant Tile_X7Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X8Y2, LUT4AB
constant Tile_X8Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000";
--X9Y2, RAM_IO
constant Tile_X9Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y3, W_IO
constant Tile_X0Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101111110010000000000000000000";
--X1Y3, LUT4AB
constant Tile_X1Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000101000000000";
--X2Y3, LUT4AB
constant Tile_X2Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X3Y3, RegFile
constant Tile_X3Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y3, LUT4AB
constant Tile_X4Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X5Y3, LUT4AB
constant Tile_X5Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X6Y3, DSP_top
constant Tile_X6Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y3, LUT4AB
constant Tile_X7Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X8Y3, LUT4AB
constant Tile_X8Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000";
--X9Y3, RAM_IO
constant Tile_X9Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y4, W_IO
constant Tile_X0Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000011101011110110000000000000000000";
--X1Y4, LUT4AB
constant Tile_X1Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000110000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001001000000000110000000000000000000000000000001000000000000";
--X2Y4, LUT4AB
constant Tile_X2Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000";
--X3Y4, RegFile
constant Tile_X3Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y4, LUT4AB
constant Tile_X4Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000";
--X5Y4, LUT4AB
constant Tile_X5Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X6Y4, DSP_bot
constant Tile_X6Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y4, LUT4AB
constant Tile_X7Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X8Y4, LUT4AB
constant Tile_X8Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X9Y4, RAM_IO
constant Tile_X9Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y5, W_IO
constant Tile_X0Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101011110111000000000000000000";
--X1Y5, LUT4AB
constant Tile_X1Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000";
--X2Y5, LUT4AB
constant Tile_X2Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X3Y5, RegFile
constant Tile_X3Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y5, LUT4AB
constant Tile_X4Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X5Y5, LUT4AB
constant Tile_X5Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X6Y5, DSP_top
constant Tile_X6Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000000000000000000000000000000000000000000000000000000000000000000";
--X7Y5, LUT4AB
constant Tile_X7Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X8Y5, LUT4AB
constant Tile_X8Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X9Y5, RAM_IO
constant Tile_X9Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y6, W_IO
constant Tile_X0Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100101110100000000000000000000";
--X1Y6, LUT4AB
constant Tile_X1Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X2Y6, LUT4AB
constant Tile_X2Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X3Y6, RegFile
constant Tile_X3Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y6, LUT4AB
constant Tile_X4Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X5Y6, LUT4AB
constant Tile_X5Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000";
--X6Y6, DSP_bot
constant Tile_X6Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y6, LUT4AB
constant Tile_X7Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X8Y6, LUT4AB
constant Tile_X8Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X9Y6, RAM_IO
constant Tile_X9Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y7, W_IO
constant Tile_X0Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000011110111110110000000000000000000";
--X1Y7, LUT4AB
constant Tile_X1Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000001000000100000000000000000000000100000000010010000000100000000010000000000000000000000000000000000000000011000000000000000000001000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000011000000000000000";
--X2Y7, LUT4AB
constant Tile_X2Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000001000000000";
--X3Y7, RegFile
constant Tile_X3Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000";
--X4Y7, LUT4AB
constant Tile_X4Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X5Y7, LUT4AB
constant Tile_X5Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000001000000000000000000000000000001011111000000000000000000000000001100101000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000100000000000000010000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000";
--X6Y7, DSP_top
constant Tile_X6Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000001101000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000";
--X7Y7, LUT4AB
constant Tile_X7Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000001000000000000000010100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000011001000000000000000000000000010000000100000000000000000000000000000000010000000000000000000000000000000000100000000000000000000000000001000000000000010000000000000000000000000000110000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000000000000000000";
--X8Y7, LUT4AB
constant Tile_X8Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000";
--X9Y7, RAM_IO
constant Tile_X9Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y8, W_IO
constant Tile_X0Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000011101011110001000000000000000000";
--X1Y8, LUT4AB
constant Tile_X1Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000001010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000100000000000000000000000000000000000010000000000000000000010000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000100000000000";
--X2Y8, LUT4AB
constant Tile_X2Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X3Y8, RegFile
constant Tile_X3Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y8, LUT4AB
constant Tile_X4Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X5Y8, LUT4AB
constant Tile_X5Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000100000000000000000000000000000111010000000000000000000000010010000000010000000100000000000000000000000000000010001000110100000010001000000100000000110000000000011101001000000000101101000000000010000000000000000101000000010011000101000000001100001000010000001000000000000000000000001000000000000110000000000100011001100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000010000000011000011000000000000000000001001100000100001001000000010000000000000000000000001000000000";
--X6Y8, DSP_bot
constant Tile_X6Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000110100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000100000000000000000011000000000000000000000000000000";
--X7Y8, LUT4AB
constant Tile_X7Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000100000000000000000000000000000000000000000000000000000000100000000000000000100000000100010010110000000000000100001000001000001100000000100110000010011010000000001000000000000000111000000000000000000100001000000000000000000000000001000000000000000000000000000001000000000001100000000001100000010001000000000000100100000000000001000010100100001000100000000000000010110000000000001100000000000010100010000001001000000000000001111000000000000100000000000001100000010000000010000000001001001100000000000010100000001000000000000100000000000000000000001111010000000000000000000000001011000100011000000000000000000100000000000000000010000";
--X8Y8, LUT4AB
constant Tile_X8Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000001000001000000000000000010001000000000000000000000000001001010010000110000001110000100000100001000110100000000010000000001100000001000000000010110100000010000000100100000000100001100001110000000000000000000000000101011010000010000000100000010010110000000000000000010100000001111000000000000000001100011100000000000100000101000000010011000000101000000000000000010010100000001001000000010000000000010000000000000000000000110001000100000000100100000000010000110000000000000000000000000010000000000010100100000011000000110100000000010010000000001011001000100010001100000000000010011101001001000000000000000000000000000001000000000000";
--X9Y8, RAM_IO
constant Tile_X9Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y9, W_IO
constant Tile_X0Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111110111000000000000000000";
--X1Y9, LUT4AB
constant Tile_X1Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000100000000000";
--X2Y9, LUT4AB
constant Tile_X2Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X3Y9, RegFile
constant Tile_X3Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000";
--X4Y9, LUT4AB
constant Tile_X4Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000010000001000000000000001000000000000000000100000100000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000110000000000000000010000000000100000010000000000000000000000000000000000000000000000000000000000000000010000000000000";
--X5Y9, LUT4AB
constant Tile_X5Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000100000000000000010100000010000010000000000000000110000000000000011000000000000000000000000000000001001000000000000100000010000000000001100010010000001000000001000101110001000001000000000010010110010101011010000000000000100000000011001001000010000000000000000001010111000000000000001100000000011000101000000000000011000000000011001101010000000000010000000000000101110000000000100000010001000010110000000000000100000000100000000000000000000000000100000000100001000000000001100000001000000100100000001000100001100100000010010000000011001001101100010001100000000000100000001001000110000000000000000000000000000000011010001";
--X6Y9, DSP_top
constant Tile_X6Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000101000000000000011010000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000011000000000000000000000000000000";
--X7Y9, LUT4AB
constant Tile_X7Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000111111000000000000001000010001100000000000000000000000100000100011001000000100010000000000000100000110000000110001100000000000000010010010000000000111010000001100100011000000000000000000000000000011010000000100000010111000000000110000110000001000001000100000000000000000000000000000000000011001010010000000000000000000010100001000010000000001000000000000100000100110010000000000000110010000001010000000000000010101011000000000000000100001000001000010000000011010000000011000101101000011110000000000000110000100000010000000000000011011001101100100001000000001000100000000001001110000100000000000000000000000000001100000";
--X8Y9, LUT4AB
constant Tile_X8Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001000000000000000000000000010001000000001000000001010101000000001000000000000000100110000000000000001101000000000000000011010000010000001000000010000000000000001100000111001000010110001010000000000000110010000100000000100000001011000100001000000000000011000000000100000011000000000000000100010011000111011000001110000011101100101000010100000000000001100000100000100000010000000101100000000000001111000000000000000000011000000000000000000000000000100011000100001000000001100100001100001011100000000001010110000101100000000010000000001010001010110101001000000000001001011101001000000000000000000000000000100000001011000010";
--X9Y9, RAM_IO
constant Tile_X9Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001010100000000000000000000000000000000000000000100000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000";
--X0Y10, W_IO
constant Tile_X0Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001101100100000000000000000000";
--X1Y10, LUT4AB
constant Tile_X1Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000";
--X2Y10, LUT4AB
constant Tile_X2Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X3Y10, RegFile
constant Tile_X3Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y10, LUT4AB
constant Tile_X4Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000100000000000000000000000000010000000110000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X5Y10, LUT4AB
constant Tile_X5Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000010001000001000000000000000000000110000010010000000000000000000000000000010000010000100000000000100010000001011000000110000000100001000000010010000000010000011000111001000000010000000000110001000000000001000011000000100000000000000100001010010110000000000101100000000001000000000000000000001000000001111000010000000001100101000001111011101010101000000000000000111000101100001000000010000000010011000000111000000000010011100000000000000100000000000010000100000001000011000000000000100000000001000000100000001000111000001100010000000000000010010001100011010000000000000000010000100001000010000000000000000000000000001000100110010";
--X6Y10, DSP_bot
constant Tile_X6Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y10, LUT4AB
constant Tile_X7Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011000000000000000011000000000000000010000000001100001011000000000000110010001001000000000000001100000000000110000000010000000011000000001010000001100010001000000100010000000000000001000001000000100000010000000000011010001001000010000001001000000010000011010000000001100001000001111101011101000000100100000000011000000011001001000000000010001100000000110100000000000010000111000000010000100000010000101000010000001000000000000001000100000001000011000000001001100011101000011000100000000100110000100100110000010000000011001011101100001000000000000000010000110010010010010000000000000000000000001000000000000";
--X8Y10, LUT4AB
constant Tile_X8Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000101000000000001100011000000000101011111000000001100110000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000001000000000000000000010000000000001100000000000000000000000000000000100110000000000000000000000000000001010100001000000000000000000000000110000100001000011000000000000001000100000000000000010000100001010000000000000000000000000000010000000000000110000010000011000100000000000000000000100000000000000000010101100000000101000000000000000000000000011011000000000000000000000000000000000011010000";
--X9Y10, RAM_IO
constant Tile_X9Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000111000111000000000000000000000000000010000000000000100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000001000000010";
--X0Y11, W_IO
constant Tile_X0Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000111101001111110000000000000000000";
--X1Y11, LUT4AB
constant Tile_X1Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000";
--X2Y11, LUT4AB
constant Tile_X2Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000";
--X3Y11, RegFile
constant Tile_X3Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000";
--X4Y11, LUT4AB
constant Tile_X4Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X5Y11, LUT4AB
constant Tile_X5Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000010000100100000000000010001000000000000000000000000100000000000000000001000000000101110000000000000100000000000000100000000001100100000000100011010000000000000000000000100010000000000000000000000000001000011000000000000000000000000000000001111000000000000000000000000000000000000000000000010000001100010011100000000000001000000010100000110000001000000001000000000000001000110000000000010100000000001000000000000000000000000010000000000000011100000000101100000000000000000000000000010101001011000000000000000000001111000000000000000000000000011000010000000000000000000001010000000000001000000000000000000000000001000011100000";
--X6Y11, DSP_top
constant Tile_X6Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y11, LUT4AB
constant Tile_X7Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000100000000101010000001010011011000000000001000010010000110000001010000100000100001100000100000000010000000001100000011000000000011010010000000000111000101000000000001000000000000000111100000000001000000000010000010110101100010101000000000110001100011100000001010011000010000010100101000011100010100001000101000100000011111011001011000000001001100010000000001100111000000010000000101010000010010000000000000100010000000100001101000000000000000110000000000001100000001001000001000011000010100000000000110100101100100010000000000001100001100111010101100000000001110000001000000011000000000000000000000110001000100100000";
--X8Y11, LUT4AB
constant Tile_X8Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000001100000010100100000110100000001000001010001000000001000010101110100010001010010100000100111001001011000000010000000000100000000000000100010010000000010100000000101001101000001101001000110100000000100000001000110001100000110000000000000001110111000101000000001100001001010011000000000000000010100001111000101010000010110100010001111101001011001000000000001000110100100000111010000000001110000110000101000011001110000010100000100000000100001000010010000100000000010010010011000000110011100000111100100000000000010010010100010000010000000011001001011100001001000000000001010011101010011000000000000000000000000111001000011010010";
--X9Y11, RAM_IO
constant Tile_X9Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000001100000000000101010100000000000000000000000001000010000000000000000100000000000000000000110000000000000001000100000000000000000011011101110101110000000000000000011000011010000000000000011111110000100100000100010000101011111110000000110010001010000000000000";
--X0Y12, W_IO
constant Tile_X0Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000000000000011111111111110000000000000000000";
--X1Y12, LUT4AB
constant Tile_X1Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X2Y12, LUT4AB
constant Tile_X2Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000010000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000010000000000000000000000000000001000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000000000000000000000000000001110011000000000000000000000000010000000000101000000000";
--X3Y12, RegFile
constant Tile_X3Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000100000000010";
--X4Y12, LUT4AB
constant Tile_X4Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011000000000000000000000000000000000000001000000000";
--X5Y12, LUT4AB
constant Tile_X5Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000001000000000001100000000000000000000110001001010000000000000000001010000100000100010100000000001100000000000000000001001000001101100000000110000000000001000000010000100110000100000000100001000001010000001000100001100000010000110000010000000000000000000110000000000000001000000001000000000000000000000001000001100000000010010000110100000000000110101000000010000000000011100000101000000011000010010100000100000001000000000000000110000000111100000000000011000000000110000000101010000000000001000000001100011100100000000000100000001100000000000000000000001001010010011001000000000001110101111010001000000000000000000000000000001001011000000";
--X6Y12, DSP_bot
constant Tile_X6Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000011000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010";
--X7Y12, LUT4AB
constant Tile_X7Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000100000000000000000000000000000000000100000000000000000000000000100000101000000000000000000000000100100100010000000000000000001000000000001000001000000000000000000110000000000000000000000100000000010000000010000000000000000000001000000000000000000100001000000000100100010010000010000000100000000010000000000100100001100000000000000000001110000000000000000000000000000000000001000";
--X8Y12, LUT4AB
constant Tile_X8Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000111001011000001000000000000000000000000000000010010101000000000000000000010000011100100100010010101000101010001001110000001010101000110001110000001000000000110100000110110001000000000000000101100010000100000001000001001010100000000001000100010000001111000110100000100101001100001000000000001101100000000000000100001000000110100000000010011100000010010000001110010000100000100000111010010001110001101001000101000011000110010101110011000001000101000000001001100010000000011000000010001000100000111011000100101000000000011000000000011110000000000010001010100000000001100000000010000100100110001100000000000000000000000001000000000000000";
--X9Y12, RAM_IO
constant Tile_X9Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000001101010000000000000001001100011011001111010000000000000000000000000100000100100001000000000001010000000000000001000111010101011111110000000000000000000000001010100010111111101111110010001001000000000101001111111110000000111000001001111100001001";
end package emulate_bitstream;
