library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package emulate_bitstream is
--X0Y1, W_IO
constant Tile_X0Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000";
--X1Y1, LUT4AB
constant Tile_X1Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100001000000000000010101010000000000111010000000001001001010100111101100111000000001000001111111101001100000000000000000000111000011110101000011000100000000100100000001000000001000000000000000100100000011001010000000000000011001010000010001001000000001111110000000000000000000000000010010100000010000000001100000001000001000010000000000000000000010000100000000000000000110100000000000010000000000000000000000000000000000000000000000000100000001000000000000000000010000000000000000001100000011000100000010000000000000100000000000000000001000011000000001000000000000001100000010000000000000000000000000000000000000000011010000";
--X2Y1, LUT4AB
constant Tile_X2Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000110000000000010101010000000111110001100000001001001010100110011100110110000001000001111110100001100000000000000000000111000011110100001010000000000000100101001100000100001000000000000111000100000000000010000000000000010000010000000000000000000001011010000000010000000000000000001110100000110000001000000000000000000000010000100000000000000000000100000000000000000000000000010100000000000000001010000000000010000000000000000000000000000000000000000000000000001000000000001000000000000011000000000010100110001100100000000000000000001000000100000000000000000000000000011011000100000010000000000000000000000000000001000000";
--X3Y1, RegFile
constant Tile_X3Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000";
--X4Y1, LUT4AB
constant Tile_X4Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000011000000000000000000000000000000111110001100000000001101111100100011010110110000000000110111100010101011100000000001000000111111001010100000000001000000100010100000000000000000000000000000101000000000000100000000010000000110001010000100000000000000000011000000000001000000000000000011110111000001100000000100000000000011000001100100001000001000000000100010000000000000000100000000100010000000000001000000000000010000000000000000000000000000000000000000010000000000000000000000000000100000000010000000011000000000001100000000000000000000100000000010001000000000000000010011000000000000000000000000000000000000000000000000000";
--X5Y1, LUT4AB
constant Tile_X5Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000110000000000011110000000100100000000000000001000001111010111011100111110000001000001101111100001111000010000000000000111000010000101000000000000000010100110000000000000000000000000000110110000000000000000000000000000111101100000100000000000000000010010000000000000000000000000001100100000010000000100000000001000101010010011000000000000000000000000000100000000000000000000000000011000000000010000000000000000100000000000000000000000000000000000000000000000010000000000000000000100000011110100000011000000000000000000010000000000001101011000000000001100000000000000000010011000100000000000000000000000000000001001000000";
--X6Y1, DSP_top
constant Tile_X6Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000";
--X7Y1, LUT4AB
constant Tile_X7Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000010000000000000000000000100100101001010000001001101111010001011100101100000001000001111111110001111000010000000000000111011000000100000000000000000000101100100000001000000000000010000000000000000100000000000100000000010001100000101000000000000001111011000000000010000000000000011110100000000000000000000000001100000000000000100000000000000000000100001000000000000110000000000100000000000000001000000000000011100000000000000000000000000000000000100000000000010000000000000000011100001011010100000000000010000000000000000000000000000000001010000000000000000000000100001100000001100000000000000000100000000000000011000000";
--X8Y1, LUT4AB
constant Tile_X8Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000001000000000000000000000000000100100110001100000001101101111010111011100110110000010000111111111100001100000000000001000000100010011110100000011000000000100000100000000000000000000001000000101110100000000000001010010000000111101000000000000000000000000010001000000000000000000000000011100101000011100000000100000000000101000010011000000000010000000000100010000000000000000100000000000011100000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000100000000010000000000000000000000010000000001010000000000010001000000000000010000001001000000000000000000000000000000001001000000000";
--X9Y1, RAM_IO
constant Tile_X9Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y2, W_IO
constant Tile_X0Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001100000000000000000000000";
--X1Y2, LUT4AB
constant Tile_X1Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100001100000000000010101010000000000111010000000000001000010100101101010111000000010000101111101011101011100000000000001000110001001010101000000000000000010110100000000000000000000000000000110000000000000000000000000000000110001010000100000000000000000011011000000001000100011000000001110110000000000000000000000001010100000000011110000000000000000000000000100100001000000000000000100101000100000001000000000000010000010000000000000000000000000000000000000000000000000000000000000000100000011010000000011000000000000000000000000000000010100000000000000000000000000000100111000100000000000000000000000000000000000000001000000";
--X2Y2, LUT4AB
constant Tile_X2Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000010101010000000111000000000000001001001010100110011100111110000001000001111110000001111000010000000000000111001100000101001000000000000100101010000000000100001000000000000101110000000001000110000000000000111101110000000000000000000000010001000000000000000000000000011100110010010000000000010000000010100000010011000000000000000000000100000110000000000000010000000000100000000000100000000000000000100000000000000000000000000000000000000000000000000000000001000000010100000000000000000001000000000000100000010010000000001000000000000001000100000000000000111010000000000000000000000000000000000000000000010000";
--X3Y2, RegFile
constant Tile_X3Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y2, LUT4AB
constant Tile_X4Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011110000000100100110001100000000000001111010111011100110110000000000110101111000001111000000000000000000111101100000100000000000000000000011000000100000000100001000000000111100000000000000100001000000000011000100000100000000000000001011110000000000000010000000000000010110100000011000000000000000000000000001100000000000000000000000100000000000000000000000000010000000010000000000000000000000000100000000000000000000000000001000000000000000000010000000000000100111100000000010100000000000000000001000000000000000000000011011000011000001000000000000000000000001000000000000000000000000000000000000000000000";
--X5Y2, LUT4AB
constant Tile_X5Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000000000000011001100000100100110001100000001000001100010111011010110110000001000001111111000001011100000000000000000111011101010100000000000000000000101000001100000000000000000000000111000000001000000000000000000000001100000001000000000000000001010010000000001000000000000000001011110100000010000000000000000000000000000000011001000010000000000100000000000001100000000000010001000000000000000010000000000010000000000000000000000000000001000000000000000000001000000000000000000000000011000000000000100011010100100000000000000000000000100001000001000000000000000100000000000100010000000000000000000000000000000011010000";
--X6Y2, DSP_bot
constant Tile_X6Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y2, LUT4AB
constant Tile_X7Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000001000110000000000010101010000100100000000000000000001001010010111011010111110000000000110111111000001011100010000000000000111101101010101000000000010000010011010000000000000100001000000000110000010000000000100001000000000110001001000100000000000000000011011000000001000000000000000001110110100001100000000000000001001100000000011100001000000000000000000100000100000000000000000000100000000100000001000000000000010000000000000000000000000000000000000100000000000000000000000000000010100001011010000000000000000000000100000000000000000000000000000000001000000000000000011011000000000000010000000000000000000000000000010000000";
--X8Y2, LUT4AB
constant Tile_X8Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001001000000000011110000000100100000000000000000000000111010001011010111110100010000101101111110001011100010000000001000110001001010101010100000010000010111110000000000000000000110000000110100010000000001000000000000000111001000000000001001000000000011110000000000000100000000000000010100000000000000001000000001100100000000011000000100010000000000000000000000000001001000000000000000000010000000000000000000001010001100000000000100000000001010000100000000100000000000000000000000100000000000000000000000000010100000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000100000";
--X9Y2, RAM_IO
constant Tile_X9Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y3, W_IO
constant Tile_X0Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001100000000000000000000000";
--X1Y3, LUT4AB
constant Tile_X1Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011110000000000111110001100000000000001111100110010000110110000000000110101110000001110110000000001000000111101101100100000000000000000100011000001100000001000000000000000101000000000000000000000010000000110001110000001000000000000000011000000000000010011000000000011110111000000000000000000000000000000000001100000000001000000000000100010000000001000110000000000100000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000001000000001010000000000000001000000000001100010010000000000011101000000010000001100000000000100000010111000000000000000000000000000000000001000000000";
--X2Y3, LUT4AB
constant Tile_X2Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011001100001000110111010000000000000000100010110001100111000000010000101110111101001111000000000010001000110010010000101000100000000000000110100000000000000000000000100000000000000001000000000000000000000001101110001000000000000000001110011000000000000000000000000011011100000000011000000010000001010000000000000100000000000000000000100001000000000000001010000000000100010110000001000000000000010100000000000000000100000000001001000100000000000010000000001100100000000000000000100000011010000100000000000010000000000000000001000000000000100000000000000011000100001010000000000000000000000000000000000000000";
--X3Y3, RegFile
constant Tile_X3Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y3, LUT4AB
constant Tile_X4Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001000000000000010101010000100100111010000000000001001010010111011100111000000000000110111111000001111000000000000000000111101100000101000000000000000100011000000001000001001000001000000101000000000001000111010000000000110001100000000100001000000000011000000110000010011010000000011110110000000000010001010000000010001000000000000000001010000000000100000001100000000000010000000100100000000000000000000000000010100000100100000000000000000000000000110000000000000000000000000000000100000000000000000000000001000000100000000010000000001000000000000010000000000000000000000011000000000000000000000000000000000000000100000000";
--X5Y3, LUT4AB
constant Tile_X5Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000010000000000010101010000000111101001010000001101001010100110011010101100000010000111111110000001011100010000000000000100001101010100000000001000000100001000000000000010000000000000000101000001000000000000000100000000110001010000000000000000000000011001000000101000000000000000011110110000000000000000100000000000011000000000110001000001000000000100001000100001000000100000000100000000000000001000000000000010010000000000000000000000000000000000000000000000000000000000010010000000000011000000000000000000000000100000000010000000000000000000000000000000000000000101101000000000001000000000000000000000000000000011100000";
--X6Y3, DSP_top
constant Tile_X6Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y3, LUT4AB
constant Tile_X7Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011110000000000000110001100000000000000111100111101010110110000010000101101111001001011100000000000001000110001101010100000000000100000100111000001100010000000001000000000101000000001000000100001000000000101101010011000000000000000000010000000000001000000000000000011011110100000011000010001000000001000000001100000001010000000000000100000000000000000000000000000000000000000000000000000000000010001000000000000001000000000001001000000000000000000000000000000100000000000000000000000001000001000111100000000000000000000100011000100001000000000000000000000000000001000010000000000000000000000000000000000000";
--X8Y3, LUT4AB
constant Tile_X8Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100001000000000000011001100000000000000000000000001100001100100001101100111110100110000111111111111001100000010000100000000100011001110101110000000000000000001110000000100010000000000000000000100100000000011000000000000000011001010000010000110000000001111110000000000000000000000000010010100000010000000010000000001000000000010000010000110000000000000100000000000001001001000000000000000000010000000000000000000001010101000000000000100000000001010000000000000000000000000000000000000100000000000000000000000000001100000000000000000000001000001000000000000000000000000100000011000000001000000000000000000000000000000000100000";
--X9Y3, RAM_IO
constant Tile_X9Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y4, W_IO
constant Tile_X0Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001100000000000000000000000";
--X1Y4, LUT4AB
constant Tile_X1Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011110000000100100101001010000001000001111010111011100101100000001000001101111100001111000010000000000000111000010000100001000000000000010100100000000000100001000000010000110000000000000000010000100000000110001100000000000000000000000011010000000000000000000000000001110100000000000010000000000001100101000000011100000000000000000000000000011000000000000010000000100000000000000001000000000000010100000100000000000000000000000000001100000000100000000000000000000100000000000010000000011000000000000100000010000000000000000000000000000000100000000000000111100000000000000000000000000000000000000000000010000";
--X2Y4, LUT4AB
constant Tile_X2Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001000000000000000000000001000110110001100000001101101111010110000000110110000010000111110111101001110110000000001000000100010011100100000000000000000100000100100000001010000000000000000101100000000100111000000010000000111001110000000001001000000000011100000000000000001000000000010010101000000000000011000000000000000000001100000000001000000000000100010000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000000001000001101000000000000000011000010000001000000010000000000001000000110010000000100000000000001011000000000000000000000000000000000000000001000000000";
--X3Y4, RegFile
constant Tile_X3Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y4, LUT4AB
constant Tile_X4Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000000000000011001100000100100000000000000001100001100010111011100111110000110000111111111000001100000010000000100000100011101110101000000000010000000001010000000000010100001000000000111110100001000010100001000000000011100000000000000110000000001010010000000010100000000000000001100110100000000001110000000000000000000000000000000010100000000000100100000000000000000000000010001000000000000000011000000000000010000100000100000000000000000000000100000000000001000000001010000000000000000010000000001100010000000000000000000000000000100011000000000000000000000001100000000000101000000000000000000000000000000000000000000";
--X5Y4, LUT4AB
constant Tile_X5Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000110100000000010101010000100100111010000000000001001010010101011100111000000000000110111101010101100000000000100000000111101001110101000000000000000010010100000000000000000000001000000110100110000000000001010000000000111001000000000000000000000000011110000000000001000000000000000010110000001000000000000000001000001000001100000100000110000000000000000010000000000000000000000000011000001000000101000000000000000000000000000000000000000001000000000000000000010000000000000000000000000011000100000011000000011111000000000000000000000000001000000010000000000000000000000000000000101000000000000000000000000000000001100000";
--X6Y4, DSP_bot
constant Tile_X6Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y4, LUT4AB
constant Tile_X7Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000111010000000000000000000000000000111110001100000000001100111100110010000110110000010000101111110000001110110000001000001000110011101100100000000010000000000111000001100000000100001000000000000000000000010000100001000000000001101110000010000000000000001110010000000000000100000000000011011111100001100000000000000001001011000000000000000000000000000000100010000000000100110000000000000010000000000000000000000000010000010000010000000000000000001000000000000100000000000000000001000000001000000000000000000000000011100000000010000000000000000000000000000000000000000000110000000000000000000000000000000000000000000010000000000";
--X8Y4, LUT4AB
constant Tile_X8Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000100000000011110000000100100110001100000001100001111010111011010110110000010000111101111100001011100000000000000000100000011010100000011000000000000000100001100000010000000000000000000000000000010010000000000000000001101000000010000000000000001110010001000000000000000000000011011100000000011000010100000001000001000000000000000010010000000000100000001000000000110100000000000010000000000000000000000000010001000100000000000000000000001001000100000000000000000000000000100000000001000100000000010000000001100000000000000000000010000001000100000001000000000000100000000011000000000000000000000000000000000000000100000";
--X9Y4, RAM_IO
constant Tile_X9Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y5, W_IO
constant Tile_X0Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010101101111000000000000000000";
--X1Y5, LUT4AB
constant Tile_X1Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000001000000000000000000000000000000000111111010000000001101101111100000011010111000000010000111111110110001011100000000000000000100011001010101000000000000000100001100100000000000000000000000000101110000000100000000000000000000111101010000000000000000000000010001000000000000000011000000011100100000001100000000000000000010100000001111000000010001000000000100001000000000000000000000000000101000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000010100000000100000000001000010000001000000000000000000000011000010011000001000000000000010000000101000000000000000000000000000001000000000000000";
--X2Y5, LUT4AB
constant Tile_X2Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011001100000000111111010000000001000001100100110011010111000000001000001111110100001011100000000000000000111010011010101000011000000000000100100000000000000000000000000000111110000001000000000000000000000011100010001000000000000000001010010000000000000000010000000001100100000000011000000100000000000111000000011000000000000000000000100000100000000000000100100010000000000000000000000000000000000001001000000000000000000000000001000000000000000000000000001000111100000000011000000000011000001100000100000010000000000000100000001000001000100000000000000000000000000000000000000000000000000000000100001010000";
--X3Y5, RegFile
constant Tile_X3Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y5, LUT4AB
constant Tile_X4Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000010101010000100100101001010000000001000010010111010000101100000010000101111111100001110110010000000001000110000011100100000011000000000100110100001100000000000000001000000101110000001001000001010000000000111101100001000100001000000000010000100000001100000000000000011100100000000000000101100000000000011000000000000001000110000000000100000000000000000000100000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000000000000011100000000000000000011000001000100100000000010000000000000000000000010000000000000000000000000100000010010000000000000000000000000000000000000";
--X5Y5, LUT4AB
constant Tile_X5Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000010000000100000000010101010000100100110001100000000001001010010101011100110110000000000110111101010101111000000000001000000111101000000100000000000000000000010100000001000000001000001000000111000000000001000011010010000000001100100000100000000000000001010010000000010000000000000000001011111000001110001000000000000000000000000000000000000010000000000110010000000000000000000000010000000000000000000010000000000010100000000100000000000000000001000000010000000000011000000000001000000001000000000100000010000010000000100000000000000000000000001110000011000000000000000010000000000000001010000000000000000000000000000000100000";
--X6Y5, DSP_top
constant Tile_X6Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y5, LUT4AB
constant Tile_X7Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000011000000000000000000000000000000111110001100000000001100111100110011100110110000010000101111110100001100000000000000001000110010011110100000011000000000000110100001000000000000000000000000000000100000000000000000000000000010000010000000000000000000000011000000000000000000000000000001110000000011100000000100000000000001000010000100000000000000000000000000000000000000000100000000100010000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000010100100000010000000000001000000000100000000100000000000011011001000000000010000000000000000000000000001000000000";
--X8Y5, LUT4AB
constant Tile_X8Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011001100000100100110001100000000000000100010001011010110110000010000101111111110001011100000000001001000110011001010100000100000000000000111100000000000000000000111000000111100000001000001001010000000000011000000001000001001000000001011110000000010000100000000000000010100000000000001001000000000100000000000000000000100010000000000100000000000000001000000000010000000000001000000010000000000001000000000100000000000000000001000000100000000000001000000000000000001100001000000000000000000011010101000000000000000000000001000001110010000000000000000000000100011000000000010000000000000000000000000000000000";
--X9Y5, RAM_IO
constant Tile_X9Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y6, W_IO
constant Tile_X0Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011101101110000000000000000000";
--X1Y6, LUT4AB
constant Tile_X1Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000001000000000000000000000000000000111111010000000000001101111100110011100111000000000000110111110000001111000000000000000000111111100000101000000000000000000011000000000001000100000000000000000110000000000100000000000000000011101110000000000000000000001110011000000000000001011000000011100110000001100000100000000001010000000000000100000001000001000000100001000100000000000000000000000100100000000001000000000000000100000000000001000000000000000000000000000000000010000000000000000000001000000000100000000100000000000000000010000000000001000011000010000000000000000000011001011000110000000000000000000000000000000000001000000";
--X2Y6, LUT4AB
constant Tile_X2Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001010000000000000000000000000111000000000000000001101111100000011100111110000000000110111000000001100000010000000000000111110001110101000000001010000010010010000000001000000000000000000110100110000000101000000000000000111001011000000001001000000000011110000000000000001000000000000010100000001100000001100000001000101000010011000000001001000000000000000100000000000000100000000000011000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000001000000000000000000000000000000011101000000000000000000000000000000000000001000011000000";
--X3Y6, RegFile
constant Tile_X3Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000";
--X4Y6, LUT4AB
constant Tile_X4Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000000000000011110000000000000110001100000000000001111100111100000110110000000000110101111101001110110000000001000000111100011100100000011000000000000010100001100010001000000000000000111110000000000000000000010000000011100110000000000000000000001010011000000010100011000000000001100101000000000001100100000000000001000000000010000001100000000000100010000000001000000100000010000010100100000000011000000000000000000000000000001000000000000000000000000000000001000000000001000000000000000000000000011000110011100000000000000000000011000000100000000000000000000000000000010000000000000000000000000000000000000000000000000";
--X5Y6, LUT4AB
constant Tile_X5Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011110000000100100101001010000001100001111010101010000101100000010000111101101010101110110010000000000000100001001100100000000010000000000000100000000010000000000001000000111100000000000001001010000000000011000100000100000000000000001011111000000001000000000000000000010110100000011000010000000000000000000000000000001010010000000000100101000000000000000000000010000000010000000000000000000000000000000000100000001000000000001000000010000000000000000000000000000011100000000110000000010000000000000100000000000000000000000011000000010001000000000000000000000001000100010000000000000000000000000000000000000";
--X6Y6, DSP_bot
constant Tile_X6Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y6, LUT4AB
constant Tile_X7Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000100000000000010101010000000111101001010000000001000010100000011100101100000110000101111110110001100000010000100001000110001001110100000100000000000000111100100000000000000000000000000111000100000100000000000000000000010000010000000000110000000001011010000000001000100000000000001110100000000001000000000000000000000000000000100001100000000000000100000000000000001000000000010100000000001000001000000000000011010000000000000000000000000000010000010000000000000000000001000000000000000011000000000001000110010100100000010000000000000100000000000010000100000000000000001000000000000010000000000000000000000000000001010000";
--X8Y6, LUT4AB
constant Tile_X8Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011001100000000111000000000000001000001100100110011100111110000001000001111110000001100000010000000000000111011101110101000000000010000100101011000000000000000000000000000101000100001000000000000000000000101101010001000000000000000000010001000000000000000000000000011011110100010000000000000000000000000000010000011000000001000000000100100000100001100000000000000000000000001000000010000000000010000000000000000000000000000001000000000000000000001000000000000000000000000011000000000000000011000000000000000000000000011000000110000010000000000000001100000010000000010000000000000000000000000000001101000000";
--X9Y6, RAM_IO
constant Tile_X9Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y7, W_IO
constant Tile_X0Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000101100010000000000000000000";
--X1Y7, LUT4AB
constant Tile_X1Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000100000000000011001100001000110110001100000000000000100010110001100110110000110000101110111101001100000000000101001000110010011110100100010000000000100110100100000100000000000000000000101000100001100000000000010000000110001010001000000110000000000011000000000000000000000000000011110101000000000000000000000000000000000001100100000100000000000000100010000000000001000000000000110000000000000001000000000000010010000000010000000000000000000010000000000000000000000000000001000000001000000000000000011000110000101000000000000000000000100100000111000000000000000000000001000000000010000000000000000000000000000000111000000";
--X2Y7, LUT4AB
constant Tile_X2Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000001000000000000000010101010000000111000000000000000001001010100000011010111110000000000110111110110001011100010000000000000111101001010101000000001000000010011110000000000000000000110000000110100000000000000000000000000000111001010000000000000000000000011110000000000000000000000000000010100000011100000000100000001100001000011100000100000101000000000000000001000000000000100000000000010001000000000101000000000001000000000000000000000000000001000100100000000000000000000001000000000000001011000000000001000000000001000000000000000000001000000000001000000000000000000010000100100000000000000000000000000000000001001001000000";
--X3Y7, RegFile
constant Tile_X3Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y7, LUT4AB
constant Tile_X4Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011110000000000000101001010000001100001111100111101100101100000110000111101111001001100000010000100000000100001101110100000000000000000000001000000000010010100001000000000111100101000000000100001000000000011000010010000001110000000001011110000000011000000000000000000010110100000000001010001000000001000000000000000001010000000000000100000000000000000000000000010001000000010001000010000000000000010000000000000001000000000001010000000000000000001000000000000000100000000000000000000000100110000000100000000000000000000000101100000001000000000000000000000000000000100000000000000000000000000000000000000000";
--X5Y7, LUT4AB
constant Tile_X5Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001000100000000000000000000100100110001100000001001101111010001011010110110000001000001111111110001011100000000001000000111011001010100000000000000000010101100100000001000000000110000000110000000010000000000000010000000110001000000101000000000000000011010000000000000000000000000001110101000000000000000000000001100100000000011000000000000000000000000010100000000000000000000000100001000000000000000000000000011000000000000000000000000000000000000100000000000000000000000000000101100001011010000000000000000000000100000000000000000000010000000000000000000000000000000000100001000001000000000000000000000000000000011100000";
--X6Y7, DSP_top
constant Tile_X6Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y7, LUT4AB
constant Tile_X7Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011110000000100100110001100000001000001111010111011100110110000101000001101111100001100000000000101000000111000011110100001011000000000100100100000000010100001000001000000101100100000000000011010010000000111001000000000000110000000000011100000000000000000000000000010010101000000000000010100000000000011000001100000000010010000000000100010000000000000000100000000010010000000000000000000000000000010000000110000001000000000001010000010000000000000000000000001000000000000000000000000010000000000011100000000010000000000010001000010010000000000000000000000000001000000000000000000000000000000000000000010000";
--X8Y7, LUT4AB
constant Tile_X8Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000010101010000000111000000000000000001000010100110011100111110000010000101111110000001100000010000100101000110001101110101000100000010000000111010000001000000001000000000000111000110000001000010000000000000001100010000000000110000000001010010000000000000100000000000001011110000000011000000000000000000000000000000011000100000000000000100000000000001001000000000010010000000000000000000000000000010011000100000000000000000000001010000100000000100000000000000000101100000000000000000000000000000010101100000010000000000010000000000100000000100000000000100000000000000000000000000000000000000000000000000010000";
--X9Y7, RAM_IO
constant Tile_X9Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y8, W_IO
constant Tile_X0Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001100000000000000000000000";
--X1Y8, LUT4AB
constant Tile_X1Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011110000000000000000000000000001100001111100101101010111110000010000111101101011101011100010000000100000100001001010101000000000110000100000110000000010000000001100000000101110000000000000000001000000000111101010000100100110000000000010000000000100100000000000000011100110100000000000110001000000000000000000000000000010100000000000100000000010000000000000000000011000000000000000001000000000000010010000000000001000000000000000100000000000000000000000000010000000000000000010000000011000001000000000000000000000000000100011001000000001000000000000000000000000000010000000000000000000000001000000000100000";
--X2Y8, LUT4AB
constant Tile_X2Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000010000000000000000000000000000100100110001100000001001101111010001011100110110100001000001111111110001111000000000001000000111011000000100010000000000000000101100000000000000000000000000000000110000000000000000000010000000011101100000000000000000000001110010001000000000000000000000011100101000001100000100010000001000000010000000100000000010000000000100010000000000000001000000000000000000011000001000000000000001100101000010000000100000000000000000000000000000000000000000001000000001000011000000000001000001000000000000000000000000000100000001000010010000000000000010101000100000010001000000000000000000000000000001000000";
--X3Y8, RegFile
constant Tile_X3Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y8, LUT4AB
constant Tile_X4Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000000000000000000000000000000111010000000001101101111100101101010111000000010000111111101011101011100000000000000000100011001010101000000000100000000000100000000000000000001100000000111100000000000010001011000000000011000010000000010000000000001011110000000100001000000000000000010110100001011000000001000000001000000001100000000000000000000000100000000000000000000000000010000000000001000000000000000000000001010000000000000000000000001000000010000000000010000000000000100000000000000000100000010100000000000010000000000000000000000101000000010000000000000001100000000000001000000000000000000000000000000000000000000";
--X5Y8, LUT4AB
constant Tile_X5Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000000000000011110000000000000101001010000001000001111100001101100101100000001000001101111111001100000010000000000000111001001110100001000000000000100101100100000010100001000000010000101000100100100000010000100000000110001010000001000000000000000011001010000000010000000000000011110100000000000000000000000000100001000010000010000000000000000000100000000000001000010000000000100010000100000000000000000000011000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000010000000100000000010000000010000011000000000000000000000000100000100000000100010000000000000000000000000000000010000";
--X6Y8, DSP_bot
constant Tile_X6Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y8, LUT4AB
constant Tile_X7Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000011000000011001100000000111101001010000001100001100100000011100101100100010000111111110110001100000010000000000000100011001110100010000001000000000001100000000100010000000000010000111000100100000000000000100000000001100010000000000000000000001010010000000010000000000000000001011100000010011001000100000000100011000010000000000000001000000000100000000000000000001100000010000000000010000000010000000000011001101000000000000100000000001000000100000000100001000000000100100000000001000000000000000000010000000000000000000000000001000000000000000000000000000000000000111000000000000000000000000000000000000000000000000";
--X8Y8, LUT4AB
constant Tile_X8Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000000000000011110000000000000000000000000001100001111100111101100111110000010000111101111101001100000010000000100000100000011110101000000000010000010000110000000000010000000000000000110110100000000010000000000000000111101010000000000110000000000010010000000000100000000000000001100100000000000000110000000001000100000010011010000010100000000000000000010100001000000000000000010000000000000000001000000000000010000000000000001000000000000010000000000000000000000000001000000000000000000000000000011000000000000100000000000000000001000001000000000000000000000000100000001000000000010000000000000000000000000001000010000";
--X9Y8, RAM_IO
constant Tile_X9Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y9, W_IO
constant Tile_X0Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000101100010000000000000000000";
--X1Y9, LUT4AB
constant Tile_X1Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011001100001000110101001010000000000000100010110000000101100000010000101110111001000000000010000010001000110011100000100000100000000000000111000000000000000000000000100000111110000001000000000000000000000011100010001000000000000000001010010000000010100100000000000001100110100000000001100000000000000100000000000010000100100000000000110100100000001001001000000010000000000010000000011001000000000010100001000000000100000000000000001000000000000001000000000000000100000000000000000000001000110111100000000000000000000000100000100000000000000000000000000000000000000010000000000000000000000000010000000000000";
--X2Y9, LUT4AB
constant Tile_X2Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000000000000011110000000000000110001100000000000000111100101101100110110000010000101101101011101100000000000000001000110001001110100000000000000000000110100001100000000000000000000000111000100001000000000000000000000001100010001100000000000000001010011000000000000000000000000001011110000010011000000000000000000000000010000011000000000000000000100000000000001100000000000010000000000100000000010000000000010001000000000000000000000000001000000000000000000001000000000000100000100000000010000000010000111000100000000000000000000011000000000100000001000000000000100000011000000010000000000000000000000000000000000000000";
--X3Y9, RegFile
constant Tile_X3Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y9, LUT4AB
constant Tile_X4Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000001000000000000011110000000100100000000000000001100001111010111011010111110000010000111101111100001011100010000000000000100000011010101000000000000000100000110000000000010000000100000000101000000000000010000000000000000110001000000001100001000000000011000000000100010000000000000011110100000010000000011000000000000000000010000000000010010000000000100000000000000000110000000000100000010000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000010100000000100000000011100000000000000000010010000000001011011000000000001100000000001100000010101001000000000000000000000000000000001000000000";
--X5Y9, LUT4AB
constant Tile_X5Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000001000000000000000000100100101001010000000001100111010001010000101100000010000101111111110001110110010000000001000110011001100100000000000000000000111100101000001000000000000000000111100000010100000000000000000000011000100000000000000000000001011110000000001000100000000000000010100000000011000000000000000000001000001100000001000000000000000100000000000000000000000000010000000010000000000000000000000001000000100000000000000000000001000000100000000000000000000000000100000000001000000000000000100110000111100000000000000000000000000100110000000000000000000000000000000110000010000000000000000000000000000000000000";
--X6Y9, DSP_top
constant Tile_X6Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y9, LUT4AB
constant Tile_X7Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000000000000011001100000000000110001100000001100001100100111101100110110000010000111111111001001111000000000001000000100011100000100100000000000000010001000000000100010100001000000000110000001100000000100001010000000101101110000000000000000000000010010000000000000000000000000001011111100000000000000000000001001100000000011010000100000000000000000010000000001101000000000000001001000000000000000000000000010100000000010000000000000000001000000000000100000000000000000001000000000000000000000000000100000001100000000000000000000000000101000000000000000000000000100000000000010000000000000000000000000000000000000000000";
--X8Y9, LUT4AB
constant Tile_X8Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000010000010000000000010101010000000000111010000000000001000010100111100000111000000010000101111111001001110110000001000001000110001101100101000000010000000000111000000000000000100001000000000111000000001000000100001000000000001100110011000000000000000001010011000000000000000011000000001011111100000011000000001000000010000000000000001000000000000000000100111000000000100000000000010001100000000000000010000000000010000000000010000000000000000001000000000000000000001000000000001000010100000011000000000000000011000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000001000011000000";
--X9Y9, RAM_IO
constant Tile_X9Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y10, W_IO
constant Tile_X0Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001001100100000000000000000000";
--X1Y10, LUT4AB
constant Tile_X1Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000010000000011000000000000000000000111111010000000000001100111100110010000111000000010000101111110100001110110000000000001000110010011100101000011000000000100110100001100000000000000000000000101000000000000000000000000000000101101110000000100001000000000010000000000000000100000000000011011100000001111000001100000000000001000000000000000000000000000000100000001000000000000100000000000010010000000000000000000000010000000000000000000000000000001001000000000000000010000000000000100011100000000000100000011000000010100000000010010000000010000011000000000000100000000000010000000000000100000000000000000000000000000000000000000";
--X2Y10, LUT4AB
constant Tile_X2Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000000000000010101010000000000101001010000000001001010100001101010101100100000000110111111111001011100010000000000000111101001010100010000000000000000011100000001000000001000000010000000000000000011000010000100000000010001010010010000000000000001111010000000000000000000000000011110100000001100000000001000001100000000000000100000000000000000000100000000000000000111000000000100000000010000001000000000000011000101100000000000100000000000000000100000000000000000000000000000000000001000000000000000000000000000100000000000000000001001000000000001000000000000001110101100001000000000000000000000000000000000001000000000";
--X3Y10, RegFile
constant Tile_X3Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y10, LUT4AB
constant Tile_X4Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000001000000000011110000000000000101001010000001100001111100111101010101100000010000111101111001001011100010000000000000100001101010100000000000100000000001000000000010000000001100010000111100000000000001000001100000000011000010000000000000000000001011110000000010000000000000000000010110110000000001010001000000100000000000000010000010000000000000100100000000001000000000000010001000000000000000010000000000000000000100000000001000000000001000000100000000000001000000010000001100000001000100000001000000110000000000000000000000000000011001100000000001000000000001100000100000000000000000000000000000000000000000000100000";
--X5Y10, LUT4AB
constant Tile_X5Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000001000000000000000011001100000000111101001010000000000001100100000011010101100100000000110111110110001011100010000000000000111111001010100010000001000000000011100000000000000000000100000100000000000001010000000000000000000001101010000010000000000000001110010000000101000000000000000011011100000001100000000100000001000001000000000000001000001000000000100000001000000000111100000000000000000010000000000000000000011000100011000000000100000000001000000010000000000000000000000000000000010000000000000000000100000100000100000000000000000000000000000000010000000000000000010000000000000000010000000000000000000000001000000000000";
--X6Y10, DSP_bot
constant Tile_X6Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y10, LUT4AB
constant Tile_X7Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000001000000011001100000000000000000000000001100001100100111101010111110000010000111111111101001011100010000000100000100010011010101000011000000000100000110000000100000000000110000000101100000000000000000000000000000111001010000000000000000000000011101000000000000000000000000010010100010000000000000100000000100111000001100010000000000000000000100000101100001000000100000000000001000100000000000000000000000000000000001000000000000000001000000100000000100000000000000000000011100000000100000000010000000000001000000000010000000000100000000000000001000000000001100000100011000000000000000000000000000000000000000000000";
--X8Y10, LUT4AB
constant Tile_X8Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000100000000000000000011110000000000000111010000000000000000111100111100000111000000010000101101111001001110110000000000001000110001101100101000000000100000000111000001100010000000001000000000000000000001000000000001000000000001101110001000000000000000001110011000000000000000011000000011011110100000000000010001000001010000000000000111000010000000000000100000000000001000000000000000000100000100000001000000000000010000000000000000001000000000001000000000000000000000000000000000000000000000000000000000000000001011100000000000000000000000000001000000000000000000000000100000000000000110000000000000000000000000000000111000000";
--X9Y10, RAM_IO
constant Tile_X9Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y11, W_IO
constant Tile_X0Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001011100101000000000000000000";
--X1Y11, LUT4AB
constant Tile_X1Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000001000000000000000011110000000100100000000000000001000001111010111010000111110000001000001101111100001110110010001000100000111000011100101000000010000000000100110000000000100000000001000000111100000000000000001010000000000011000100000000000000000000001011110000000010000000000000000000010101000000000001000000000000000000000001100000000000010000000000100010000000000000000000000010000000000000000000010000000000000000000000010100000000000000001000000000000000000001000000000001000000000000000100000000011100010000011000000010000000000000111100100000010001100000000000000000000001010000000000000000000000000000001000000000000";
--X2Y11, LUT4AB
constant Tile_X2Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011110000000000111101001010000000000000111100000011010101100100010000101101110110001011100010000000001000110001001010100010000000000000010111100000000000000000000000010000110000000001000000000000100000000110001010001001000000000000000011010000000001010000000000000001110100000000000000000000000001100000000000000000001000000000000000000000000000000000111000000000100000000010000010100000000000011000100000000000000100000000000000000100000000100000000000000000000000000000000100000000000000001000001100000000000000000000010000000000001001000000000000000000100011000010010000000000000000000000000000000000000";
--X3Y11, RegFile
constant Tile_X3Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y11, LUT4AB
constant Tile_X4Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000001000000000011110000000000000101001010000001100001111100101101010101100000010000111101101011101011100010000000000000100001001010100000000000100000010000100000000010000000001110000000110000001000000000000001000000000110001010000001000000000000000011010000000001010000000000000001110110100000000000000001000001101000000000000000101000100000000000000100000000000000110000000000100000000000000000101000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000100000000011000000000000100000000000000000010111000000000000001000000000000100000100101000000010000000000000000000000000000000100000";
--X5Y11, LUT4AB
constant Tile_X5Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000100000000000010101010001000110000000000000001101001010010110001100111110000010000111110111101001100000010000010100000100000011110101000001000010000010000110000000000000000000000100000110110100000000000000000000000000111101010000000000110000000000010010000000000000000000000000001100100000010000000100000000001000100000010011000000000000000000000000000100000000000001000000000000001000010000000000000000000000010001000000000000100000000000000000000000000000000000000000010000000000000011100000000010000000100000000001100000000000001001000000000010001000000000000000000001001000000000000000000000000000000000001001000000";
--X6Y11, DSP_top
constant Tile_X6Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y11, LUT4AB
constant Tile_X7Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000011110000000000111000000000000001100001111100110011010111110000010000111101110000001011100010000000000000100001101010101000000000010000000001010000000000010100001000000000111110010000000010100001000000000011100010000000000000000000001010010000000010100000000000000001100110100000000001110000000000000000000000000000001010101000000000100000000000000000000000000010000000000000000000011000000000000000000000000000000000000000000000001000000000000001000000001000001100000000000000000000001000010000000000000000000000000000000001110000000001000000000001100000000000001000000000000000000000000000000000000000000";
--X8Y11, LUT4AB
constant Tile_X8Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000010000000000000000011001100000000111110001100000000000001100100100011100110110000100000110111100010101100000000000100000000111111001110100000000001000000000010100001100000000000000000000000111000100000000000001010000000000001100010000000010110000000001010010000000010001000000000000001011110000001111001000100000000000011000000000000000000001000000000100000000000000000000100000010000010000000000000010000000000010011000000100000000000000000001000000010000000000001000000000000000000000000000000000000010000010010100100000000000000000000000000110000011000000000000000010000000000000000010000000000000000000000000000000000000";
--X9Y11, RAM_IO
constant Tile_X9Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y12, W_IO
constant Tile_X0Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y12, LUT4AB
constant Tile_X1Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000111000000000011110000000100100111010000000001000001111010101011010111000000001000001101101010101011100000000000000000111001001010101000000000000000000100100000000010000000000111000000000100000000000000001010000000000011001000000000000000000000001111111000000000001000011000000010010110001000000000010000000001110000000001100100000010010000000000100001000000000000000000000000000100000100000001000000000000000000000100100000001000000000001000000110000000100000000000000000000000000000011000000000010000000000001000000000000000000000000011000000010000000000000000000101100000000000000000000000000000000000000000001100000";
--X2Y12, LUT4AB
constant Tile_X2Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000010000000000000000000000000001000110101001010000001101101111010110001100101100000010000111110111101001100000010000010000000100010011110100000011000000000100000100000000000000000000000110000101110100000000000000000100000000111101010000000000000000000000010000000000000100000000000000011100100000011100000100100000000100011000011100000000000100000000000100000001000000000000100000000000000000000000000001000000000000000000000000000000100000000000000000100000000100000000000000000000000100000000100000000011000000000011000000000000000000001000000000000000000000000000000010000101100000000000000000000000000000000001000000000000";
--X3Y12, RegFile
constant Tile_X3Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000";
--X4Y12, LUT4AB
constant Tile_X4Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000110000000000000000000000000000000000000000000000001100111100111101010111110000010000101111111101001011100010000000101000110010011010101000000000100000010110110000000001000000001000000000110000000001000100000001000000000110001010001000000000000000000011010000000001000001000000000001110100100000000000000001000001000100000000011100001001000000000000000100000000000000000000000000100001000000000001000000000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000011000000000000100000010000000000001100000000000001000100000000000000001001000000010010000000000000000000000000010000000000";
--X5Y12, LUT4AB
constant Tile_X5Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000010000000000000000000000000000101001010000001101101111100111100000101100000010000111111111101001110110010001000000000100010011100100000011010100000000000100000000001000000001000000000000100000000000100000001000000000011001110000000001000000000001111110000000001000001000000000010010101100000000000000101000001000011000000000100001001000000000000100110000010000000000100000000001000000000000001000000000000000000000000010000000000000000001000000000000000000000000000000001000000000000000100000000010000000000000100000000000000000001001000000000000001000000000000000001000011000000010000000000000000000000000001011000000";
--X6Y12, DSP_bot
constant Tile_X6Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X7Y12, LUT4AB
constant Tile_X7Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000010000000000000000000000000111101001010000000001100111100000011100101100100010000101111110110001100000010000000001000110011001110100010000001000000010111100000000000000000000000010000110000100001000000000000100000000101101010001000000000000000000010010000000000000000000000000001011100000001100000000100000001100001000010000001100000101000000000000000001000000100001100000000000010000010000000111000000000011000111100000000000100000000001000000100000000000001000000000000000000000000000000000000001000011000000000000000000000000000000000011000000000000000000000000000100100000000000000000000000000000000001000111000000";
--X8Y12, LUT4AB
constant Tile_X8Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000001000110101001010000000000001000010100001010101100000000000110000101011101011100010000010000000111101001010100000000000000000000010100000000000001000000100100000000000000000000000000000000000000010000010000101000000000000000011000000000001010011000000000001110010000000000000000000000000000000000000000000001001000000000000000000000000000000111000000000100000000010000000000000000000010000100000100000000100000000000000000000000000000000000000000000000011100000000010000000010000000000000100000000000000000011000000000000010000000000000000100000000000000000010100000000000000000000000000000000000";
--X9Y12, RAM_IO
constant Tile_X9Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
end package emulate_bitstream;
